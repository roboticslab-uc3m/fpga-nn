module perceptron (
	input wire [3:0] a,
	input wire [3:0] b,
	output wire [3:0] res	
);

	assign res = a + b;

endmodule
